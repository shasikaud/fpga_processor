// module top_layer_tb();

//     reg start_sig;
//     reg [15:0] dram_in_sig;
//     reg [15:0] iram_in_sig;
//     wire [15:0] data_out_sig;
//     wire [15:0] addr_out_sig;
//     wire mem_write_sig;


// top_layer top_layer_dut
// (
// 	.start(start_sig) ,	// input  start_sig
// 	.dram_in(dram_in_sig) ,	// input [15:0] dram_in_sig
// 	.iram_in(iram_in_sig) ,	// input [15:0] iram_in_sig
// 	.data_out(data_out_sig) ,	// output [15:0] data_out_sig
// 	.addr_out(addr_out_sig) ,	// output [15:0] addr_out_sig
// 	.mem_write(mem_write_sig) 	// output [1:0] mem_write_sig
// );

// always
// 		begin
// 			#5 clock = 1;
// 			#5 clock = 0;
// 		end
		