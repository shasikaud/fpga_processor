`timescale 1ns / 1ps

module rom_vlog_mif 
#(
    parameter ADDR_WIDTH = 9,
    parameter DATA_WIDTH = 16
)
(
    input                       clk_i,
    input                     read_en,
    input                     write_en,
    input      [DATA_WIDTH-1:0]   data,
    input      [ADDR_WIDTH-1:0] addr_i,
    output reg [DATA_WIDTH-1:0] data_o
);


reg [DATA_WIDTH-1:0] mem[0:2**ADDR_WIDTH-1];

initial begin
    $readmemh("mem_init_vlog.mif", mem); 
end


always @(posedge clk_i)
begin
if (read_en == 1)begin
     data_o <= mem[addr_i];
end

if (write_en == 1)begin
     mem[addr_i] <= data;
end
   end
    
endmodule
